module CRC #(
	parameter	DATA_WIDTH = 32,
	parameter	CRC_WIDTH = 3,
	parameter	COUNTER_WIDTH = $clog2(DATA_WIDTH),
	parameter	LSB_DATA_WIDTH = DATA_WIDTH - CRC_WIDTH,
	parameter	POLYNOMIAL = 3'h3
)(
	//input	
	input								clk,
	input								reset_n,
	//control = 0, Lay gia tri luu vao thanh ghi
	//control = 1, Bat dau tinh toan
	input								control,
	input								enable,
	input		[DATA_WIDTH - 1 : 0]	data_in,
	//output
	output		[DATA_WIDTH - 1 : 0]	result,
	output	reg							done
);
	reg	[LSB_DATA_WIDTH - 1 : 0]		lsb_data_reg;
	reg	[COUNTER_WIDTH - 1 : 0]			count = 0;
	reg	[CRC_WIDTH - 1 : 0]				polynomial = POLYNOMIAL;
	reg									status;

	reg	[CRC_WIDTH - 1 : 0]				crc_result;
	wire								clear_count;
	
	//Tinh toan trang thai hien tai cua mach
	always @(posedge clk, negedge reset_n) begin
		if(~reset_n) 
			status <= 1'b0;
		else if(clear_count) 
			status <= 1'b0;
		else if(~control & enable)
			status <= 1'b1;
	end
	
	// Luu cac bit lSB vao thanh ghi result khi control = 0
	// Bat dau dich cac bit LSB khi control = 1
	always @(posedge clk) begin
		if(~control & enable)
			lsb_data_reg <= data_in[LSB_DATA_WIDTH - 1 : 0];
		else if (status & control) 
			lsb_data_reg <= lsb_data_reg << 1'b1;
		else
			lsb_data_reg <= lsb_data_reg;
	end
	
	// Bien count se dem so chu ky can de tinh CRC
	// So chu ky can dung de tinh toan CRC = so bit Data truyen vao (DATA_WIDTH)
	assign	clear_count = count == (DATA_WIDTH - 1); 
	
	always @(posedge clk, negedge reset_n) begin
		if(~reset_n)
			count <= {COUNTER_WIDTH{1'b0}};
		else if(clear_count)
			count <= {COUNTER_WIDTH{1'b0}};
		else if(status & control)
			count <= count + 1'b1;
		else
			count <= count;
	end
	
	//Sau khi dem duoc DATA_WIDTH chu ky thi se disable status = 0. Ngung tinh toan
	//Luc nay du lieu tinh toan da co the doc tu master
	always @(posedge clk, negedge reset_n) begin
		if(~reset_n)
			done <= 1'b0;
		else if(~status & control)
			done <= 1'b1;
		else 
			done <= done;
	end
	
	//Khoi tinh toan CRC o day
	always@ (posedge clk, negedge reset_n) begin
		if(~reset_n)
			crc_result <= {CRC_WIDTH{1'b0}};
		else if(~control & enable)
			//Load MSB Data tu datain vao thanh ghi  chua ket qua tinh toan CRC
			crc_result <= data_in[DATA_WIDTH - 1 : DATA_WIDTH - CRC_WIDTH];
		else if(status & control) begin
			if(crc_result[CRC_WIDTH - 1]) 
				crc_result <= {crc_result[CRC_WIDTH - 2 : 0], lsb_data_reg[LSB_DATA_WIDTH - 1]} ^ polynomial;
			else
				crc_result <= {crc_result[CRC_WIDTH - 2 : 0], lsb_data_reg[LSB_DATA_WIDTH - 1]};
		end else
			crc_result <= crc_result;
	end
	
	assign	result = done ? {{(DATA_WIDTH - CRC_WIDTH){1'b0}},crc_result} : {DATA_WIDTH{1'b0}};
	
	
	
endmodule